`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.05.2024 08:23:52
// Design Name: 
// Module Name: adder_32bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_32bit
#(
    parameter ADDER_WIDTH = 32, 
    parameter BLOCK_SIZE = 8
    )
    (
    input wire [ADDER_WIDTH-1:0] iA, iB,
    input wire iCarry,
    output wire [ADDER_WIDTH-1:0] oSum,
    output wire oCarry   
    );
    
     wire [ADDER_WIDTH/BLOCK_SIZE - 2 : 0] carry; // carry array generated by every block other than first and last because they are Cin and Cout
     assign num_of_blocks = ADDER_WIDTH / BLOCK_SIZE;
    
      genvar i;
    generate
    
      for (i = 0; i < ADDER_WIDTH/BLOCK_SIZE; i = i + 1) 
      begin : blocks
        if(i == 0)
            CLA_first 
            #( .ADDER_WIDTH(BLOCK_SIZE) ) firstBlock
            (
            .iA(iA[BLOCK_SIZE-1:0]),
            .iB(iB[BLOCK_SIZE-1:0]),
            .iCarry(iCarry),
            .oSum(oSum[BLOCK_SIZE-1:0]),
            .oCarry(carry[0]));
        else if(i != 0 & i == ADDER_WIDTH/BLOCK_SIZE - 1)
            CLA_inter 
            #( .ADDER_WIDTH(BLOCK_SIZE))  lastBlock
            (
              .iA(iA[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),
              .iB(iB[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),
              .iCarry(carry[i-1]),
              .oSum(oSum[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),          
              .oCarry(oCarry)   
            );
        else
            CLA_inter 
            #( .ADDER_WIDTH(BLOCK_SIZE)) inter 
            (
              .iA(iA[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),
              .iB(iB[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),
              .iCarry(carry[i-1]),
              .oSum(oSum[BLOCK_SIZE*i+BLOCK_SIZE-1:BLOCK_SIZE*i]),          
              .oCarry(carry[i])   
            );
      end
       endgenerate
    
    
    
    
endmodule
